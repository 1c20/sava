#this is comment
define version = "1" #in-line comment
define name = "sava"
define list = | 3,2,1 |


print("program started")


loop %list %i:
    print(%i + "~~~")
    print("-")

print("exit without errors")
